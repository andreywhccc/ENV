`define SVT_MST_IF_CONNECT(PATH,SVT_IF_INST,PORT_ID)\
    assign ``PATH``araddr                           = ``SVT_IF_INST``[``PORT_ID``].araddr   ;\
    assign ``PATH``arburst                          = ``SVT_IF_INST``[``PORT_ID``].arburst  ;\
    assign ``PATH``arcache                          = ``SVT_IF_INST``[``PORT_ID``].arcache  ;\
    assign ``PATH``arid                             = ``SVT_IF_INST``[``PORT_ID``].arid     ;\
    assign ``PATH``arlen                            = ``SVT_IF_INST``[``PORT_ID``].arlen    ;\
    assign ``PATH``arlock                           = ``SVT_IF_INST``[``PORT_ID``].arlock   ;\
    assign ``PATH``arprot                           = ``SVT_IF_INST``[``PORT_ID``].arprot   ;\
    assign ``PATH``arsize                           = ``SVT_IF_INST``[``PORT_ID``].arsize   ;\
    assign ``PATH``arvalid                          = ``SVT_IF_INST``[``PORT_ID``].arvalid  ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arready     = ``PATH``arready                       ;\
    assign ``PATH``awaddr                           = ``SVT_IF_INST``[``PORT_ID``].awaddr   ;\
    assign ``PATH``awburst                          = ``SVT_IF_INST``[``PORT_ID``].awburst  ;\
    assign ``PATH``awcache                          = ``SVT_IF_INST``[``PORT_ID``].awcache  ;\
    assign ``PATH``awid                             = ``SVT_IF_INST``[``PORT_ID``].awid     ;\
    assign ``PATH``awlen                            = ``SVT_IF_INST``[``PORT_ID``].awlen    ;\
    assign ``PATH``awlock                           = ``SVT_IF_INST``[``PORT_ID``].awlock   ;\
    assign ``PATH``awprot                           = ``SVT_IF_INST``[``PORT_ID``].awprot   ;\
    assign ``PATH``awsize                           = ``SVT_IF_INST``[``PORT_ID``].awsize   ;\
    assign ``PATH``awvalid                          = ``SVT_IF_INST``[``PORT_ID``].awvalid  ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awready     = ``PATH``awready                       ;\
    assign ``PATH``wdata                            = ``SVT_IF_INST``[``PORT_ID``].wdata    ;\
    assign ``PATH``wlast                            = ``SVT_IF_INST``[``PORT_ID``].wlast    ;\
    assign ``PATH``wstrb                            = ``SVT_IF_INST``[``PORT_ID``].wstrb    ;\
    assign ``PATH``wvalid                           = ``SVT_IF_INST``[``PORT_ID``].wvalid   ;\
    assign ``SVT_IF_INST``[``PORT_ID``].wready      = ``PATH``wready                        ;\
    assign ``PATH``bready                           = ``SVT_IF_INST``[``PORT_ID``].bready   ;\
    assign ``SVT_IF_INST``[``PORT_ID``].bid         = ``PATH``bid                           ;\
    assign ``SVT_IF_INST``[``PORT_ID``].bresp       = ``PATH``bresp                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].bvalid      = ``PATH``bvalid                        ;\
    assign ``PATH``rready                           = ``SVT_IF_INST``[``PORT_ID``].rready   ;\
    assign ``SVT_IF_INST``[``PORT_ID``].rdata       = ``PATH``rdata                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].rid         = ``PATH``rid                           ;\
    assign ``SVT_IF_INST``[``PORT_ID``].rlast       = ``PATH``rlast                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].rresp       = ``PATH``rresp                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].rvalid      = ``PATH``rvalid                        ;\


`define SVT_SLV_IF_CONNECT(PATH,SVT_IF_INST,PORT_ID)\
    assign ``SVT_IF_INST``[``PORT_ID``].araddr      = ``PATH``araddr                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arburst     = ``PATH``arburst                       ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arcache     = ``PATH``arcache                       ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arid        = ``PATH``arid                          ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arlen       = ``PATH``arlen                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arlock      = ``PATH``arlock                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arprot      = ``PATH``arprot                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arsize      = ``PATH``arsize                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arvalid     = ``PATH``arvalid                       ;\
    assign ``PATH``arready                          = ``SVT_IF_INST``[``PORT_ID``].arready  ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awaddr      = ``PATH``awaddr                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awburst     = ``PATH``awburst                       ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awcache     = ``PATH``awcache                       ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awid        = ``PATH``awid                          ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awlen       = ``PATH``awlen                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awlock      = ``PATH``awlock                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awprot      = ``PATH``awprot                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awsize      = ``PATH``awsize                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awvalid     = ``PATH``awvalid                       ;\
    assign ``PATH``awready                          = ``SVT_IF_INST``[``PORT_ID``].awready  ;\
    assign ``SVT_IF_INST``[``PORT_ID``].wdata       = ``PATH``wdata                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].wlast       = ``PATH``wlast                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].wstrb       = ``PATH``wstrb                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].wvalid      = ``PATH``wvalid                        ;\
    assign ``PATH``wready                           = ``SVT_IF_INST``[``PORT_ID``].wready   ;\
    assign ``PATH``bid                              = ``SVT_IF_INST``[``PORT_ID``].bid      ;\
    assign ``PATH``bresp                            = ``SVT_IF_INST``[``PORT_ID``].bresp    ;\
    assign ``PATH``bvalid                           = ``SVT_IF_INST``[``PORT_ID``].bvalid   ;\
    assign ``SVT_IF_INST``[``PORT_ID``].bready      = ``PATH``bready                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].rready      = ``PATH``rready                        ;\
    assign ``PATH``rdata                            = ``SVT_IF_INST``[``PORT_ID``].rdata    ;\
    assign ``PATH``rid                              = ``SVT_IF_INST``[``PORT_ID``].rid      ;\
    assign ``PATH``rlast                            = ``SVT_IF_INST``[``PORT_ID``].rlast    ;\
    assign ``PATH``rresp                            = ``SVT_IF_INST``[``PORT_ID``].rresp    ;\
    assign ``PATH``rvalid                           = ``SVT_IF_INST``[``PORT_ID``].rvalid   ;\


`define SVT_MON_IF_CONNECT(PATH,SVT_IF_INST,PORT_ID)\
    assign ``SVT_IF_INST``[``PORT_ID``].araddr      = ``PATH``araddr                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arburst     = ``PATH``arburst                       ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arcache     = ``PATH``arcache                       ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arid        = ``PATH``arid                          ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arlen       = ``PATH``arlen                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arlock      = ``PATH``arlock                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arprot      = ``PATH``arprot                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arsize      = ``PATH``arsize                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arvalid     = ``PATH``arvalid                       ;\
    assign ``SVT_IF_INST``[``PORT_ID``].arready     = ``PATH``arready                       ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awaddr      = ``PATH``awaddr                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awburst     = ``PATH``awburst                       ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awcache     = ``PATH``awcache                       ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awid        = ``PATH``awid                          ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awlen       = ``PATH``awlen                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awlock      = ``PATH``awlock                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awprot      = ``PATH``awprot                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awsize      = ``PATH``awsize                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awvalid     = ``PATH``awvalid                       ;\
    assign ``SVT_IF_INST``[``PORT_ID``].awready     = ``PATH``awready                       ;\
    assign ``SVT_IF_INST``[``PORT_ID``].wdata       = ``PATH``wdata                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].wlast       = ``PATH``wlast                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].wstrb       = ``PATH``wstrb                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].wvalid      = ``PATH``wvalid                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].wready      = ``PATH``wready                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].bid         = ``PATH``bid                           ;\
    assign ``SVT_IF_INST``[``PORT_ID``].bresp       = ``PATH``bresp                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].bvalid      = ``PATH``bvalid                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].bready      = ``PATH``bready                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].rready      = ``PATH``rready                        ;\
    assign ``SVT_IF_INST``[``PORT_ID``].rdata       = ``PATH``rdata                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].rid         = ``PATH``rid                           ;\
    assign ``SVT_IF_INST``[``PORT_ID``].rlast       = ``PATH``rlast                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].rresp       = ``PATH``rresp                         ;\
    assign ``SVT_IF_INST``[``PORT_ID``].rvalid      = ``PATH``rvalid                        ;\
